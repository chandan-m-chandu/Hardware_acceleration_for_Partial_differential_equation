
module element_tb();
logic CLK; logic R; logic [15:0]Wx; logic [15:0]Wy; logic [15:0]W;
logic [15:0]bi[4:0][4:0];
logic [15:0]uij[4:0][4:0];
PEarray uut( CLK, R, Wx, Wy,W, bi, uij);
initial
begin
CLK=0;R=1;Wx=1;Wy=1;W=1;
bi=&#39;{&#39;{0,0,0,0,0},&#39;{0,0,0,0,0},&#39;{0,0,0,0,0},&#39;{0,0,0,0,0},&#39;{0,0,0,0,0}};
uij=&#39;{&#39;{0,0,0,0,0},&#39;{0,0,0,0,0},&#39;{0,0,0,0,0},&#39;{0,0,0,0,0},&#39;{0,0,0,0,0}};
#10;R=0; bi =&#39;{&#39;{1,1,1,1,1},&#39;{1,1,1,1,1},&#39;{1,1,1,1,1},&#39;{1,1,1,1,1},&#39;{1,1,1,1,1}};
#10 CLK=1;#10 CLK=0;
#10 CLK=1;#10 CLK=0;
#10 CLK=1;#10 CLK=0;
#10 CLK=1;#10 CLK=0;
#10 CLK=1;#10 CLK=0;

#10 CLK=1;#10 CLK=0;
#10 CLK=1;#10 CLK=0;
#10 CLK=1;#10 CLK=0;
#10 CLK=1;#10 CLK=0;
#10 CLK=1;#10 CLK=0;
#10 CLK=1;#10 CLK=0;

$finish;
end
endmodule
